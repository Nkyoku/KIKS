library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

library work;
use work.misc_pkg.all;
use work.openMSP430_pkg.all;
use work.BusTest_pkg.all;


entity TestBenchOMSP is
end TestBenchOMSP;



architecture Simulation of TestBenchOMSP is
	
	signal clk_sys		: std_logic;
	
	signal reset		: std_logic;
	
	signal interval		: std_logic;
	
	signal mem_en		: std_logic := '0';
	signal mem_wr		: std_logic := '0';
	signal mem_wait		: std_logic;
	signal mem_addr		: std_logic_vector(15 downto 0) := X"0000";
	signal mem_din		: std_logic_vector(15 downto 0) := X"0000";
	signal mem_dout		: std_logic_vector(15 downto 0);

	subtype ROM_BYTE is std_logic_vector(15 downto 0);
	type ROM is array (0 to 8191) of ROM_BYTE;
	constant PROM : ROM := (
			X"0A12", X"0912", X"0943", X"0A43", X"1B43", X"0F93", X"0424", X"094D", X"0D4C", X"0C43", X"0D3C", X"0C5C", X"0D6D", X"0969", X"098E", X"0428",
			X"1CD3", X"0B5B", X"F82B", X"033C", X"095E", X"0B5B", X"F42B", X"1B43", X"0C5C", X"0D6D", X"0969", X"0A6A", X"098E", X"0A7F", X"0428", X"1CD3",
			X"0B5B", X"F62B", X"043C", X"095E", X"0A6F", X"0B5B", X"F12B", X"0E49", X"0F4A", X"3941", X"3A41", X"3041", X"0A12", X"0912", X"3F40", X"60C1",
			X"3F93", X"1224", X"3D40", X"60C1", X"0C3C", X"8F12", X"2A53", X"123C", X"3C4D", X"0A4D", X"0E49", X"B012", X"12C1", X"0A59", X"0D4A", X"1D53",
			X"1DC3", X"394D", X"0993", X"F423", X"3F40", X"FFFF", X"3F93", X"0524", X"3A40", X"FFFF", X"2F4A", X"0F93", X"E823", X"3040", X"2EC1", X"3140",
			X"0080", X"B240", X"44C1", X"4A40", X"B240", X"44C1", X"4C40", X"B012", X"3CC1", X"0C93", X"0224", X"B012", X"58C0", X"0C43", X"B012", X"EAC0",
			X"B012", X"40C1", X"0A12", X"0A43", X"0B43", X"12C3", X"0D10", X"0C10", X"0228", X"0A5E", X"0B6F", X"0E5E", X"0F6F", X"0D93", X"F623", X"0C93",
			X"F423", X"0C4A", X"0D4B", X"3A41", X"3041", X"8243", X"4200", X"B240", X"0180", X"2000", X"F240", X"1000", X"0000", X"32D2", X"FF3F", X"0E43",
			X"12C3", X"0C10", X"0128", X"0E5D", X"0D5D", X"0C93", X"F923", X"0C4E", X"3041", X"0F4C", X"0E93", X"0524", X"1F53", X"FF4D", X"FFFF", X"1E83",
			X"FB23", X"3041", X"3441", X"3541", X"3641", X"3741", X"3841", X"3941", X"3A41", X"3041", X"F240", X"1000", X"0000", X"0013", X"1C43", X"3041",
			X"0343", X"FF3F", X"3041", X"2530", X"386C", X"5800", X"2025", X"3032", X"5800", X"2025", X"3038", X"4C58", X"0000", X"2025", X"3034", X"5800",
			X"0200", X"4840", X"0100", X"0200", X"5840", X"0000", X"0100", X"3A40", X"FF00", X"0100", X"5640", X"0000", X"0000", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF",
			X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"34C1", X"9EC0"
		);
	
	

begin
	
	
	OMSP : OMSPWrapper
		generic map(
			PBUS_BASE_ADDRESS	=> X"1000"
		)
		port map(
			CLK_SYS1		=> clk_sys,
			CLK_SYS2		=> clk_sys,
			RESET			=> reset,
			OMSP_RESET		=> open,
			TICK_SYNC_IN	=> '0',
			TICK_CNT_OUT	=> open,
			NMI_IN			=> interval,
			IRQ_IN			=> "00000000000000",
			IRQ_ACC			=> open,
			PBUS_EN			=> mem_en,
			PBUS_WR			=> mem_wr,
			PBUS_WAIT		=> mem_wait,
			PBUS_ADDR		=> mem_addr,
			PBUS_DATA_IN	=> mem_din,
			PBUS_DATA_OUT	=> mem_dout,
			XBUS_EN			=> open,
			XBUS_WR			=> open,
			XBUS_ADDR		=> open,
			XBUS_DATA_IN	=> X"0000",
			XBUS_DATA_OUT	=> open,
			XDMA_EN1		=> '0',
			XDMA_EN2		=> '0',
			XDMA_WR			=> '0',
			XDMA_ADDR1		=> X"000",
			XDMA_ADDR2		=> X"000",
			XDMA_DATA_IN	=> X"00000000",
			XDMA_DATA_OUT1	=> open,
			XDMA_DATA_OUT2	=> open
		);
	
	
	
	-- クロック生成(50MHz)
	CLK1_process : process begin
		clk_sys <= '1';
		wait for 10.000 ns;
		clk_sys <= '0';
		wait for 10.000 ns;
	end process;
	
	-- Interval生成
	Interval_process : process begin
		interval <= '0';
		wait for 10 us;
		wait until rising_edge(clk_sys);
		interval <= '1';
		wait until rising_edge(clk_sys);
	end process;
	
	
	
	
	-- データ生成
	-- Signal_process : process begin
		
		
		
		
		
		-- wait for 500 us;
		-- assert (false) report "Simulation End" severity failure;
		-- wait;
	-- end process;
	
	-- バス信号生成
	Bus_process : process begin
		-- リセット
		reset		<= '1';
		wait for 100 ns;
		reset		<= '0';
		wait for 100 ns;
		
		wait for 1 us;
		
		-- バスアクセス
		BusWrite(CLK_SYS, mem_en, mem_wr, mem_addr, mem_din, X"1000", X"0002");
		wait for 1 us;
		for cnt in 0 to 8191 loop
			BusWrite(CLK_SYS, mem_en, mem_wr, mem_addr, mem_din, X"1001", PROM(cnt)(15 downto 8) & PROM(cnt)(7 downto 0));
		end loop;
		wait for 1 us;
		BusWrite(CLK_SYS, mem_en, mem_wr, mem_addr, mem_din, X"1000", X"0003");
		
		wait for 100 us;
		assert (false) report "Simulation End" severity failure;
		wait;
	end process;
	
end;
